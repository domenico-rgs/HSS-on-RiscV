// File             : log_param.vh
// Author           : D. Ragusa
// Creation Date    : 11.01.24
// Last Modified    : 11.01.24
// Version          : 1.0
// Abstract         : Constants and parameters for the Log Module

`define COEFF_FILE "data_file/log_coeff.hex"
`define PIPE_NREG 3
`define DECIMAL_BITS 12