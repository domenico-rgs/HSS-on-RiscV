// File             : butterworth_const.vh
// Author           : D. Ragusa
// Creation Date    : 11.01.24
// Last Modified    : 11.01.24
// Version          : 1.0
// Abstract         : Constants and parameters for the Butterworth Low-pass filter

`define COEFF_FILE "data_file/butter_coeff.hex"
`define DECIMAL_BITS 12
`define N_COEFF 3
