// File             : exp_param.vh
// Author           : D. Ragusa
// Creation Date    : 11.01.24
// Last Modified    : 11.01.24
// Version          : 1.0
// Abstract         : Constants and parameters for the Exp Module

`define COEFF_FILE "mem_files/exp_coeff.mem"
`define PIPE_NREG 3
`define ONE 16'd4096
`define DECIMAL_BITS 12