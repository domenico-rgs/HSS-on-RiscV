// File             : homo_config.vh
// Author           : D. Ragusa
// Creation Date    : 11.01.24
// Last Modified    : 11.01.24
// Version          : 1.0
// Abstract         : Constants and parameters for the Homomorphic Chain Module

`define LOG_N_STAGES 2
`define ONE 16'h1000
`define EXP_N_STAGES 2